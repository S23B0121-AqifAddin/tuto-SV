import streamlit as st 

  st.set_page_config(
    page_title="Scientific Visualization"
  )

  st.header("Scientific Visualization", divider="grey")
